class master_seq_r extends uvm_sequencer #(master_seq_i);

    `uvm_component_utils(master_seq_r)

    function new(string name="master_seq_r",uvm_component parent=null);
        super.new(name,parent);
    endfunction

    


endclass