package elv_pkg;
 `include "master_seq.sv"
    

endpackage 