class slave_seq_r extends uvm_sequence;

    `uvm_component_utils(slave_seq_r)
    function new(string name="slave_seq_r",uvm_component parent=null);
    super.new(name,parent);
    endfunction


endclass